module Strip (
    input logic [31:0] in,
    input logic signal,
    output logic [31:0] out
);
    assign out = in;
endmodule