module Extend (
    input logic [31:0] in,
    input logic signal,
    input logic [31:0] out
);
    assign out = in;
endmodule